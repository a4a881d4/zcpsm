library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity crc8_blkrom is
	port(
		clk		:	in std_logic;
		addr	:	in	std_logic_vector(7 downto 0);
		dout	:	out	std_logic_vector(31 downto 0)
		);
end entity;

architecture behavior of crc8_blkrom is
	
	type array256x32 is array(0 to 255) of std_logic_vector(31 downto 0);
	constant data_array	:	array256x32	:=	(
	"00000000000000000000000000000000",
	"00000100110000010001110110110111",
	"00001001100000100011101101101110",
	"00001101010000110010011011011001",
	"00010011000001000111011011011100",
	"00010111110001010110101101101011",
	"00011010100001100100110110110010",
	"00011110010001110101000000000101",
	"00100110000010001110110110111000",
	"00100010110010011111000000001111",
	"00101111100010101101011011010110",
	"00101011010010111100101101100001",
	"00110101000011001001101101100100",
	"00110001110011011000011011010011",
	"00111100100011101010000000001010",
	"00111000010011111011110110111101",
	"01001100000100011101101101110000",
	"01001000110100001100011011000111",
	"01000101100100111110000000011110",
	"01000001010100101111110110101001",
	"01011111000101011010110110101100",
	"01011011110101001011000000011011",
	"01010110100101111001011011000010",
	"01010010010101101000101101110101",
	"01101010000110010011011011001000",
	"01101110110110000010101101111111",
	"01100011100110110000110110100110",
	"01100111010110100001000000010001",
	"01111001000111010100000000010100",
	"01111101110111000101110110100011",
	"01110000100111110111101101111010",
	"01110100010111100110011011001101",
	"10011000001000111011011011100000",
	"10011100111000101010101101010111",
	"10010001101000011000110110001110",
	"10010101011000001001000000111001",
	"10001011001001111100000000111100",
	"10001111111001101101110110001011",
	"10000010101001011111101101010010",
	"10000110011001001110011011100101",
	"10111110001010110101101101011000",
	"10111010111010100100011011101111",
	"10110111101010010110000000110110",
	"10110011011010000111110110000001",
	"10101101001011110010110110000100",
	"10101001111011100011000000110011",
	"10100100101011010001011011101010",
	"10100000011011000000101101011101",
	"11010100001100100110110110010000",
	"11010000111100110111000000100111",
	"11011101101100000101011011111110",
	"11011001011100010100101101001001",
	"11000111001101100001101101001100",
	"11000011111101110000011011111011",
	"11001110101101000010000000100010",
	"11001010011101010011110110010101",
	"11110010001110101000000000101000",
	"11110110111110111001110110011111",
	"11111011101110001011101101000110",
	"11111111011110011010011011110001",
	"11100001001111101111011011110100",
	"11100101111111111110101101000011",
	"11101000101111001100110110011010",
	"11101100011111011101000000101101",
	"00110100100001100111000001110111",
	"00110000010001110110110111000000",
	"00111101000001000100101100011001",
	"00111001110001010101011010101110",
	"00100111100000100000011010101011",
	"00100011010000110001101100011100",
	"00101110000000000011110111000101",
	"00101010110000010010000001110010",
	"00010010100011101001110111001111",
	"00010110010011111000000001111000",
	"00011011000011001010011010100001",
	"00011111110011011011101100010110",
	"00000001100010101110101100010011",
	"00000101010010111111011010100100",
	"00001000000010001101000001111101",
	"00001100110010011100110111001010",
	"01111000100101111010101100000111",
	"01111100010101101011011010110000",
	"01110001000101011001000001101001",
	"01110101110101001000110111011110",
	"01101011100100111101110111011011",
	"01101111010100101100000001101100",
	"01100010000100011110011010110101",
	"01100110110100001111101100000010",
	"01011110100111110100011010111111",
	"01011010010111100101101100001000",
	"01010111000111010111110111010001",
	"01010011110111000110000001100110",
	"01001101100110110011000001100011",
	"01001001010110100010110111010100",
	"01000100000110010000101100001101",
	"01000000110110000001011010111010",
	"10101100101001011100011010010111",
	"10101000011001001101101100100000",
	"10100101001001111111110111111001",
	"10100001111001101110000001001110",
	"10111111101000011011000001001011",
	"10111011011000001010110111111100",
	"10110110001000111000101100100101",
	"10110010111000101001011010010010",
	"10001010101011010010101100101111",
	"10001110011011000011011010011000",
	"10000011001011110001000001000001",
	"10000111111011100000110111110110",
	"10011001101010010101110111110011",
	"10011101011010000100000001000100",
	"10010000001010110110011010011101",
	"10010100111010100111101100101010",
	"11100000101101000001110111100111",
	"11100100011101010000000001010000",
	"11101001001101100010011010001001",
	"11101101111101110011101100111110",
	"11110011101100000110101100111011",
	"11110111011100010111011010001100",
	"11111010001100100101000001010101",
	"11111110111100110100110111100010",
	"11000110101111001111000001011111",
	"11000010011111011110110111101000",
	"11001111001111101100101100110001",
	"11001011111111111101011010000110",
	"11010101101110001000011010000011",
	"11010001011110011001101100110100",
	"11011100001110101011110111101101",
	"11011000111110111010000001011010",
	"01101001000011001110000011101110",
	"01101101110011011111110101011001",
	"01100000100011101101101110000000",
	"01100100010011111100011000110111",
	"01111010000010001001011000110010",
	"01111110110010011000101110000101",
	"01110011100010101010110101011100",
	"01110111010010111011000011101011",
	"01001111000001000000110101010110",
	"01001011110001010001000011100001",
	"01000110100001100011011000111000",
	"01000010010001110010101110001111",
	"01011100000000000111101110001010",
	"01011000110000010110011000111101",
	"01010101100000100100000011100100",
	"01010001010000110101110101010011",
	"00100101000111010011101110011110",
	"00100001110111000010011000101001",
	"00101100100111110000000011110000",
	"00101000010111100001110101000111",
	"00110110000110010100110101000010",
	"00110010110110000101000011110101",
	"00111111100110110111011000101100",
	"00111011010110100110101110011011",
	"00000011000101011101011000100110",
	"00000111110101001100101110010001",
	"00001010100101111110110101001000",
	"00001110010101101111000011111111",
	"00010000000100011010000011111010",
	"00010100110100001011110101001101",
	"00011001100100111001101110010100",
	"00011101010100101000011000100011",
	"11110001001011110101011000001110",
	"11110101111011100100101110111001",
	"11111000101011010110110101100000",
	"11111100011011000111000011010111",
	"11100010001010110010000011010010",
	"11100110111010100011110101100101",
	"11101011101010010001101110111100",
	"11101111011010000000011000001011",
	"11010111001001111011101110110110",
	"11010011111001101010011000000001",
	"11011110101001011000000011011000",
	"11011010011001001001110101101111",
	"11000100001000111100110101101010",
	"11000000111000101101000011011101",
	"11001101101000011111011000000100",
	"11001001011000001110101110110011",
	"10111101001111101000110101111110",
	"10111001111111111001000011001001",
	"10110100101111001011011000010000",
	"10110000011111011010101110100111",
	"10101110001110101111101110100010",
	"10101010111110111110011000010101",
	"10100111101110001100000011001100",
	"10100011011110011101110101111011",
	"10011011001101100110000011000110",
	"10011111111101110111110101110001",
	"10010010101101000101101110101000",
	"10010110011101010100011000011111",
	"10001000001100100001011000011010",
	"10001100111100110000101110101101",
	"10000001101100000010110101110100",
	"10000101011100010011000011000011",
	"01011101100010101001000010011001",
	"01011001010010111000110100101110",
	"01010100000010001010101111110111",
	"01010000110010011011011001000000",
	"01001110100011101110011001000101",
	"01001010010011111111101111110010",
	"01000111000011001101110100101011",
	"01000011110011011100000010011100",
	"01111011100000100111110100100001",
	"01111111010000110110000010010110",
	"01110010000000000100011001001111",
	"01110110110000010101101111111000",
	"01101000100001100000101111111101",
	"01101100010001110001011001001010",
	"01100001000001000011000010010011",
	"01100101110001010010110100100100",
	"00010001100110110100101111101001",
	"00010101010110100101011001011110",
	"00011000000110010111000010000111",
	"00011100110110000110110100110000",
	"00000010100111110011110100110101",
	"00000110010111100010000010000010",
	"00001011000111010000011001011011",
	"00001111110111000001101111101100",
	"00110111100100111010011001010001",
	"00110011010100101011101111100110",
	"00111110000100011001110100111111",
	"00111010110100001000000010001000",
	"00100100100101111101000010001101",
	"00100000010101101100110100111010",
	"00101101000101011110101111100011",
	"00101001110101001111011001010100",
	"11000101101010010010011001111001",
	"11000001011010000011101111001110",
	"11001100001010110001110100010111",
	"11001000111010100000000010100000",
	"11010110101011010101000010100101",
	"11010010011011000100110100010010",
	"11011111001011110110101111001011",
	"11011011111011100111011001111100",
	"11100011101000011100101111000001",
	"11100111011000001101011001110110",
	"11101010001000111111000010101111",
	"11101110111000101110110100011000",
	"11110000101001011011110100011101",
	"11110100011001001010000010101010",
	"11111001001001111000011001110011",
	"11111101111001101001101111000100",
	"10001001101110001111110100001001",
	"10001101011110011110000010111110",
	"10000000001110101100011001100111",
	"10000100111110111101101111010000",
	"10011010101111001000101111010101",
	"10011110011111011001011001100010",
	"10010011001111101011000010111011",
	"10010111111111111010110100001100",
	"10101111101100000001000010110001",
	"10101011011100010000110100000110",
	"10100110001100100010101111011111",
	"10100010111100110011011001101000",
	"10111100101101000110011001101101",
	"10111000011101010111101111011010",
	"10110101001101100101110100000011",
	"10110001111101110100000010110100");
	
begin
	
	process( clk )
	begin
		if rising_edge( clk ) then
			dout <= data_array(conv_integer(addr));	
		end if;
	end process;
end behavior;
