library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library unisim;
use unisim.vcomponents.all;
entity test is
    Port (
			addra: IN std_logic_VECTOR(9 downto 0);
			addrb: IN std_logic_VECTOR(9 downto 0);
			clka: IN std_logic;
			clkb: IN std_logic;
			dina: IN std_logic_VECTOR(15 downto 0);
			douta: OUT std_logic_VECTOR(15 downto 0);
			doutb: OUT std_logic_VECTOR(15 downto 0);
			wea: IN std_logic);
end test;
architecture low_level_definition of test is
attribute INIT_00 : string;
attribute INIT_01 : string;
attribute INIT_02 : string;
attribute INIT_03 : string;
attribute INIT_04 : string;
attribute INIT_05 : string;
attribute INIT_06 : string;
attribute INIT_07 : string;
attribute INIT_08 : string;
attribute INIT_09 : string;
attribute INIT_0A : string;
attribute INIT_0B : string;
attribute INIT_0C : string;
attribute INIT_0D : string;
attribute INIT_0E : string;
attribute INIT_0F : string;
attribute INIT_00 of ram_0 : label is  "88006301800F4301940E6001C02063018009430194086001C0200F0002010300";
attribute INIT_01 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_02 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_03 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_04 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_05 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_06 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_07 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_08 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_09 of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_0A of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_0B of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_0C of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_0D of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_0E of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_0F of ram_0 : label is  "0000000000000000000000000000000000000000000000000000000000000000";
begin
  ram_0: RAMB4_s16_s16
  generic map (
               INIT_00 => X"88006301800F4301940E6001C02063018009430194086001C0200F0002010300",
               INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
               INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
               )
  port map(
  	DIA    => dina,
        DIB    => "0000000000000000",
        ENA    => '1',
        ENB    => '1',
        WEA    => wea,
        WEB    => '0',
        RSTA   => '0',
        RSTB   => '0',
        CLKA   => clka,
        CLKB   => clkb,
        ADDRA  => addra( 7 downto 0),
        ADDRB  => addrb( 7 downto 0),
        DOA    => douta,
        DOB    => doutb
        );
end low_level_definition;
