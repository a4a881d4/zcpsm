library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package Eth_TestSig_Cfg is 
	
	signal g_Test_EthRec_CRCFlag					: std_logic; -- ethrx_input; DFE_TR 
	
end package;
